
module soc_system (
	clk_clk,
	hdmi_clk,
	reset_reset_n,
	pll_locked_export);	

	input		clk_clk;
	output		hdmi_clk;
	input		reset_reset_n;
	output		pll_locked_export;
endmodule
